`timescale 1ns / 1ps

/*
decode.sv:

  This module decodes dots and dashes into 
*/